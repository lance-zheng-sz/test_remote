module test();



endmodule
